library IEEE; 
use IEEE.STD_LOGIC_1164.ALL; 
use IEEE.NUMERIC_STD.ALL;

entity CRC8 is 
port( Clk: in std_logic; 
        reset : in std_logic; --active high reset
        size_data : in unsigned(15 downto 0);  --the size of input stream in bits.
        Data_in : in std_logic; --serial input
        crc_out : out unsigned(7 downto 0); --8 bit crc checksum
        crc_ready : out std_logic --high when the calculation is done.
        ); 
end CRC8; 

architecture Behavioral of CRC8 is 

signal count : unsigned(15 downto 0) := (others => '0');
signal crc_temp : unsigned(7 downto 0) := (others => '0');

begin

process(Clk,reset)
begin
    if(reset = '1') then
        crc_temp <= (others => '0');
        count <= (others => '0');
        crc_ready <= '0';
    elsif(rising_edge(Clk)) then
    --crc calculation in the next four lines.
        crc_temp(0) <= Data_in xor crc_temp(7);
        crc_temp(1) <= crc_temp(0) xor crc_temp(7);
        crc_temp(2) <= crc_temp(1) xor crc_temp(7);
        crc_temp(7 downto 3) <= crc_temp(6 downto 2);
        
        count <= count + 1; --keeps track of the number of rounds
        if(count = size_data + 7) then --check when to finish the calculations
            count <= (others => '0');
            crc_ready <= '1';
        end if; 
    end if; 
end process;    

crc_out <= crc_temp;

end Behavioral;