counter_inst : counter PORT MAP (
		clk_en	 => clk_en_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
